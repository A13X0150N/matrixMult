// matrix_load.sv

import mm_defs::*;

module matrix_load (
	input clk,    // Clock
	input rst     // Synchronous reset active high
);

	import matrix_pkg::*;


endmodule : matrix_load
