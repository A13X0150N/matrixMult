// mpu_adder.sv
// ----------------------------------------------------------------------------
//   Author: Alex Olson
//     Date: June 2019
//
// Desciption:
// ----------------------------------------------------------------------------
// Method to add two matrices from registers together and place the result into
// a register.

import global_defs::*;

module mpu_adder
(
	input clk,    // Clock
	input rst     // Synchronous reset active low
	
);



endmodule