// mpu_load_store_tb.sv

import global_defs::*;

module mpu_load_store_tb;

    import mpu_pkg::*;

    mpu_bfm mpu_bfm();

    mpu_register_file matrix_register_file (
        // Control signals
        .clk                    (mpu_bfm.clk),
        .rst                    (mpu_bfm.rst),
        .reg_load_en_in         (mpu_bfm.reg_load_en),
        .reg_store_en_in        (mpu_bfm.reg_store_en),

        // To MPU load
        .reg_load_addr_in       (mpu_bfm.reg_load_addr),
        .reg_i_load_loc_in      (mpu_bfm.reg_i_load_loc),
        .reg_j_load_loc_in      (mpu_bfm.reg_j_load_loc),
        .reg_load_element_in    (mpu_bfm.reg_load_element),     
        .reg_m_size_in          (mpu_bfm.reg_m_size),
        .reg_n_size_in          (mpu_bfm.reg_n_size),

        // To MPU store
        .reg_store_addr_in      (mpu_bfm.reg_store_addr),
        .reg_i_store_loc_in     (mpu_bfm.reg_i_store_loc),
        .reg_j_store_loc_in     (mpu_bfm.reg_j_store_loc),
        .reg_store_element_out  (mpu_bfm.reg_store_element),
        .reg_store_complete_out (mpu_bfm.reg_store_complete)
    );

    mpu_load load_dut (
        // Control signals
        .clk                    (mpu_bfm.clk),
        .rst                    (mpu_bfm.rst),
        .load_en_in             (mpu_bfm.load_en),

        // To memory
        .mem_element_in         (mpu_bfm.mem_load_element),
        .mem_m_size_in          (mpu_bfm.mem_load_m_size),
        .mem_n_size_in          (mpu_bfm.mem_load_n_size),
        .mem_load_addr_in       (mpu_bfm.mem_load_addr),
        .mem_load_error_out     (mpu_bfm.mem_load_error),
        .mem_load_ack_out       (mpu_bfm.mem_load_ack),

        // To matrix register file
        .reg_load_en_out        (mpu_bfm.reg_load_en),
        .reg_load_addr_out      (mpu_bfm.reg_load_addr),
        .reg_load_element_out   (mpu_bfm.reg_load_element),
        .reg_i_load_loc_out     (mpu_bfm.reg_i_load_loc),
        .reg_j_load_loc_out     (mpu_bfm.reg_j_load_loc),
        .reg_m_size_out         (mpu_bfm.reg_m_size),
        .reg_n_size_out         (mpu_bfm.reg_n_size)

    );

    mpu_store store_dut (
        // Control signals
        .clk                    (mpu_bfm.clk),
        .rst                    (mpu_bfm.rst),
        .store_en_in            (mpu_bfm.store_en),

        // To matrix register file
        .reg_element_in         (mpu_bfm.reg_store_element),
        .reg_i_store_loc_in     (mpu_bfm.reg_i_store_loc),
        .reg_j_store_loc_in     (mpu_bfm.reg_j_store_loc),
        .reg_store_complete_in  (mpu_bfm.reg_store_complete),

        // To memory
        .mem_store_en_out       (mpu_bfm.mem_store_en),
        .mem_store_element_out  (mpu_bfm.mem_store_element),
        .mem_m_size_out         (mpu_bfm.mem_store_m_size),
        .mem_n_size_out         (mpu_bfm.mem_store_n_size)
    );

    // Test variables
    mpu_operation_t op;
    logic [FP-1:0] in_matrix [M*N];
    logic [MBITS:0] in_m;
    logic [NBITS:0] in_n;
    logic [MATRIX_REG_SIZE-1:0] matrix_addr1, matrix_addr2;

    initial begin
        mpu_bfm.reset_mpu();
        op = NOP;
        in_m = 2;
        in_n = 2;
        matrix_addr1 = 0;
        matrix_addr2 = 1;
        mpu_bfm.reg_store_addr = '0;
        foreach(in_matrix[i]) in_matrix[i] = '0;
        mpu_bfm.send_op(op, in_matrix, in_m, in_n, matrix_addr1, matrix_addr2);
        op = LOAD;
        in_matrix[0] = 32'h3f800000;        // 1.0
        in_matrix[1] = 32'h424951ec;        // 50.33
        in_matrix[2] = 32'hc0200000;        // -2.5
        in_matrix[3] = 32'h3e000000;        // 0.125
        mpu_bfm.send_op(op, in_matrix, in_m, in_n, matrix_addr1, matrix_addr2);

        @(posedge mpu_bfm.clk);
        $display("\n\tTEST MATRIX LOAD\n\t%f\t%f\n\t%f\t%f\n", 
                    $bitstoshortreal(mpu_bfm.reg_element_out[0][0]),
                    $bitstoshortreal(mpu_bfm.reg_element_out[0][1]),
                    $bitstoshortreal(mpu_bfm.reg_element_out[1][0]),
                    $bitstoshortreal(mpu_bfm.reg_element_out[1][1]));
        
        /* 
        $display("\n\tTEST MATRIX LOAD\n\t%f\t%f\n\t%f\t%f\n", 
                    $bitstoshortreal(matrix_register_file.matrix_register_array[0][0][0]),
                    $bitstoshortreal(matrix_register_file.matrix_register_array[0][0][1]),
                    $bitstoshortreal(matrix_register_file.matrix_register_array[0][1][0]),
                    $bitstoshortreal(matrix_register_file.matrix_register_array[0][1][1]));
        */
    end


endmodule : mpu_load_store_tb
