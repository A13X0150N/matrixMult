// mpu_store.sv
// register file --> external source

import global_defs::*;

module mpu_store
(
	input clk,		// Clock
	input rst		// Synchronous reset active high
);

	import mpu_pkg::*;




endmodule : mpu_store
