// matrix_fetch.sv


