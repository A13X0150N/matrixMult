// mpu_load.sv

import mm_defs::*;

module mpu_load (
	input clk,    // Clock
	input rst     // Synchronous reset active high
);

	import mpu_pkg::*;


endmodule : mpu_load
