// mpu_store.sv

import mm_defs::*;

module mpu_store (
	input clk,		// Clock
	input rst		// Synchronous reset active high
);

	import mpu_pkg::*;




endmodule : mpu_store
