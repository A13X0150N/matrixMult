// mpu_controller_tb.sv

import global_defs::*;
import mpu_data_types::*;

module mpu_controller_tb;
    import testbench_utilities::*;


endmodule : mpu_controller_tb
