// mpu_controller.sv
// ----------------------------------------------------------------------------
//   Author: Alex Olson
//     Date: June 2019
//
// Desciption:
// ----------------------------------------------------------------------------
// Controller for interfacing with memory with functional units

module mpu_controller 
(
    // Control signals
    input clk,    // Clock
    input rst,    // Synchronous reset active low


);

    









    

endmodule : mpu_controller
