// matrix_store.sv

import mm_defs::*;

module matrix_store (
	input clk,		// Clock
	input rst		// Synchronous reset active high
);

	import matrix_pkg::*;




endmodule : matrix_store
