// matrix_send.sv


