// mpu_adder.sv

import global_defs::*;

module mpu_adder
(
	input clk,    // Clock
	input rst     // Synchronous reset active low
	
);



endmodule