// matrix_send_tb.sv



