// matrix_fetch_tb.sv


