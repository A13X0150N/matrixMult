// mm_pkg.sv

package mm_pkg;
	
	typedef enum logic {FALSE, TRUE} bool;

endpackage : mm_pkg

